module util

struct BBox {
	x int
	y int
	u int
	v int
}

// pub fn (b BBox) to_tex_coords(width int, height int) (f32, f32, f32, f32) {

// }
