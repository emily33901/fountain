module main

const (
	test_chars = [
		`㈀`,
		`㈁`,
		`㈂`,
		`㈃`,
		`㈄`,
		`㈅`,
		`㈆`,
		`㈇`,
		`㈈`,
		`㈉`,
		`㈊`,
		`㈋`,
		`㈌`,
		`㈍`,
		`㈎`,
		`㈏`,
		`㈐`,
		`㈑`,
		`㈒`,
		`㈓`,
		`㈔`,
		`㈕`,
		`㈖`,
		`㈗`,
		`㈘`,
		`㈙`,
		`㈚`,
		`㈛`,
		`㈜`,
		`㈠`,
		`㈡`,
		`㈢`,
		`㈣`,
		`㈤`,
		`㈥`,
		`㈦`,
		`㈧`,
		`㈨`,
		`㈩`,
		`㈪`,
		`㈫`,
		`㈬`,
		`㈭`,
		`㈮`,
		`㈯`,
		`㈰`,
		`㈱`,
		`㈲`,
		`㈳`,
		`㈴`,
		`㈵`,
		`㈶`,
		`㈷`,
		`㈸`,
		`㈹`,
		`㈺`,
		`㈻`,
		`㈼`,
		`㈽`,
		`㈾`,
		`㈿`,
		`㉀`,
		`㉁`,
		`㉂`,
		`㉃`,
		`㉠`,
		`㉡`,
		`㉢`,
		`㉣`,
		`㉤`,
		`㉥`,
		`㉦`,
		`㉧`,
		`㉨`,
		`㉩`,
		`㉪`,
		`㉫`,
		`㉬`,
		`㉭`,
		`㉮`,
		`㉯`,
		`㉰`,
		`㉱`,
		`㉲`,
		`㉳`,
		`㉴`,
		`㉵`,
		`㉶`,
		`㉷`,
		`㉸`,
		`㉹`,
		`㉺`,
		`㉻`,
		`㉿`,
		`㊀`,
		`㊁`,
		`㊂`,
		`㊃`,
		`㊄`,
		`㊅`,
		`㊆`,
		`㊇`,
		`㊈`,
		`㊉`,
		`㊊`,
		`㊋`,
		`㊌`,
		`㊍`,
		`㊎`,
		`㊏`,
		`㊐`,
		`㊑`,
		`㊒`,
		`㊓`,
		`㊔`,
		`㊕`,
		`㊖`,
		`㊗`,
		`㊘`,
		`㊙`,
		`㊚`,
		`㊛`,
		`㊜`,
		`㊝`,
		`㊞`,
		`㊟`,
		`㊠`,
		`㊡`,
  `Ё`,  `Ђ`,  `Ѓ`,  `Є`,  `Ѕ`,  `І`,  `Ї`,  `Ј`,  `Љ`,  `Њ`,  `Ћ`,  `Ќ`,  `Ў`,  `Џ`,  `А`,  `Б`,  `В`,  `Г`,  `Д`,  `Е`,  `Ж`,  `З`,  `И`,  `Й`,  `К`,  `Л`,  `М`,  `Н`,  `О`,  `П`,  `Р`,  `С`,  `Т`,  `У`,  `Ф`,  `Х`,  `Ц`,  `Ч`,  `Ш`,  `Щ`,  `Ъ`,  `Ы`,  `Ь`,  `Э`,  `Ю`,  `Я`,  `а`,  `б`,  `в`,  `г`,  `д`,  `е`,  `ж`,  `з`,  `и`,  `й`,  `к`,  `л`,  `м`,  `н`,  `о`,  `п`,  `р`,  `с`,  `т`,  `у`,  `ф`,  `х`,  `ц`,  `ч`,  `ш`,  `щ`,  `ъ`,  `ы`,  `ь`,  `э`,  `ю`,  `я`,  `ё`,  `ђ`,  `ѓ`,  `є`,  `ѕ`,  `і`,  `ї`,  `ј`,  `љ`,  `њ`,  `ћ`,  `ќ`,  `ў`,  `џ`,  `Ѡ`,  `ѡ`,  `Ѣ`,  `ѣ`,  `Ѥ`,  `ѥ`,  `Ѧ`,  `ѧ`,  `Ѩ`,  `ѩ`,  `Ѫ`,  `ѫ`,  `Ѭ`,  `ѭ`,  `Ѯ`,  `ѯ`,  `Ѱ`,  `ѱ`,  `Ѳ`,  `ѳ`,  `Ѵ`,  `ѵ`,  `Ѷ`,  `ѷ`,  `Ѹ`,  `ѹ`,  `Ѻ`,  `ѻ`,  `Ѽ`,  `ѽ`,  `Ѿ`,  `ѿ`,  `Ҁ`,  `ҁ`,  `҂`
  `Ⴀ`,  `Ⴁ`,  `Ⴂ`,  `Ⴃ`,  `Ⴄ`,  `Ⴅ`,  `Ⴆ`,  `Ⴇ`,  `Ⴈ`,  `Ⴉ`,  `Ⴊ`,  `Ⴋ`,  `Ⴌ`,  `Ⴍ`,  `Ⴎ`,  `Ⴏ`,  `Ⴐ`,  `Ⴑ`,  `Ⴒ`,  `Ⴓ`,  `Ⴔ`,  `Ⴕ`,  `Ⴖ`,  `Ⴗ`,  `Ⴘ`,  `Ⴙ`,  `Ⴚ`,  `Ⴛ`,  `Ⴜ`,  `Ⴝ`,  `Ⴞ`,  `Ⴟ`,  `Ⴠ`,  `Ⴡ`,  `Ⴢ`,  `Ⴣ`,  `Ⴤ`,  `Ⴥ`,  `ა`,  `ბ`,  `გ`,  `დ`,  `ე`,  `ვ`,  `ზ`,  `თ`,  `ი`,  `კ`,  `ლ`,  `მ`,  `ნ`,  `ო`,  `პ`,  `ჟ`,  `რ`,  `ს`,  `ტ`,  `უ`,  `ფ`,  `ქ`,  `ღ`,  `ყ`,  `შ`,  `ჩ`,  `ც`,  `ძ`,  `წ`,  `ჭ`,  `ხ`,  `ჯ`,  `ჰ`,  `ჱ`,  `ჲ`,  `ჳ`,  `ჴ`,  `ჵ`,  `ჶ`,  `჻`
  `☀`,  `☁`,  `☂`,  `☃`,  `☄`,  `★`,  `☆`,  `☇`,  `☈`,  `☉`,  `☊`,  `☋`,  `☌`,  `☍`,  `☎`,  `☏`,  `☐`,  `☑`,  `☒`,  `☓`,  `☚`,  `☛`,  `☜`,  `☝`,  `☞`,  `☟`,  `☠`,  `☡`,  `☢`,  `☣`,  `☤`,  `☥`,  `☦`,  `☧`,  `☨`,  `☩`,  `☪`,  `☫`,  `☬`,  `☭`,  `☮`,  `☯`,  `☰`,  `☱`,  `☲`,  `☳`,  `☴`,  `☵`,  `☶`,  `☷`,  `☸`,  `☹`,  `☺`,  `☻`,  `☼`,  `☽`,  `☾`,  `☿`,  `♀`,  `♁`,  `♂`,  `♃`,  `♄`,  `♅`,  `♆`,  `♇`,  `♈`,  `♉`,  `♊`,  `♋`,  `♌`,  `♍`,  `♎`,  `♏`,  `♐`,  `♑`,  `♒`,  `♓`,  `♔`,  `♕`,  `♖`,  `♗`,  `♘`,  `♙`,  `♚`,  `♛`,  `♜`,  `♝`,  `♞`,  `♟`,  `♠`,  `♡`,  `♢`,  `♣`,  `♤`,  `♥`,  `♦`,  `♧`,  `♨`,  `♩`,  `♪`,  `♫`,  `♬`,  `♭`,  `♮`,  `♯`
  `一`,  `丁`,  `丂`,  `七`,  `丄`,  `丅`,  `丆`,  `万`,  `丈`,  `三`,  `上`,  `下`,  `丌`,  `不`,  `与`,  `丏`,  `丐`,  `丑`,  `丒`,  `专`,  `且`,  `丕`,  `世`,  `丗`,  `丘`,  `丙`,  `业`,  `丛`,  `东`,  `丝`,  `丞`,  `丟`,  `丠`,  `両`,  `丢`,  `丣`,  `两`,  `严`,  `並`,  `丧`,  `丨`,  `丩`,  `个`,  `丫`,  `丬`,  `中`,  `丮`,  `丯`,  `丰`,  `丱`,  `串`,  `丳`,  `临`,  `丵`,  `丶`,  `丷`,  `丸`,  `丹`,  `为`,  `主`,  `丼`,  `丽`,  `举`,  `丿`,  `乀`,  `乁`,  `乂`,  `乃`,  `乄`,  `久`,  `乆`,  `乇`,  `么`,  `义`,  `乊`,  `之`,  `乌`,  `乍`,  `乎`,  `乏`,  `乐`,  `乑`,  `乒`,  `乓`,  `乔`,  `乕`,  `乖`,  `乗`,  `乘`,  `乙`,  `乚`,  `乛`,  `乜`,  `九`,  `乞`,  `也`,  `习`,  `乡`,  `乢`,  `乣`,  `乤`,  `乥`,  `书`,  `乧`,  `乨`,  `乩`,  `乪`,  `乫`,  `乬`,  `乭`,  `乮`,  `乯`,  `买`,  `乱`,  `乲`,  `乳`,  `乴`,  `乵`,  `乶`,  `乷`,  `乸`,  `乹`,  `乺`,  `乻`,  `乼`,  `乽`,  `乾`,  `乿`
  `가`,  `각`,  `갂`,  `갃`,  `간`,  `갅`,  `갆`,  `갇`,  `갈`,  `갉`,  `갊`,  `갋`,  `갌`,  `갍`,  `갎`,  `갏`,  `감`,  `갑`,  `값`,  `갓`,  `갔`,  `강`,  `갖`,  `갗`,  `갘`,  `같`,  `갚`,  `갛`,  `개`,  `객`,  `갞`,  `갟`,  `갠`,  `갡`,  `갢`,  `갣`,  `갤`,  `갥`,  `갦`,  `갧`,  `갨`,  `갩`,  `갪`,  `갫`,  `갬`,  `갭`,  `갮`,  `갯`,  `갰`,  `갱`,  `갲`,  `갳`,  `갴`,  `갵`,  `갶`,  `갷`,  `갸`,  `갹`,  `갺`,  `갻`,  `갼`,  `갽`,  `갾`,  `갿`,  `걀`,  `걁`,  `걂`,  `걃`,  `걄`,  `걅`,  `걆`,  `걇`,  `걈`,  `걉`,  `걊`,  `걋`,  `걌`,  `걍`,  `걎`,  `걏`,  `걐`,  `걑`,  `걒`,  `걓`,  `걔`,  `걕`,  `걖`,  `걗`,  `걘`,  `걙`,  `걚`,  `걛`,  `걜`,  `걝`,  `걞`,  `걟`,  `걠`,  `걡`,  `걢`,  `걣`,  `걤`,  `걥`,  `걦`,  `걧`,  `걨`,  `걩`,  `걪`,  `걫`,  `걬`,  `걭`,  `걮`,  `걯`,  `거`,  `걱`,  `걲`,  `걳`,  `건`,  `걵`,  `걶`,  `걷`,  `걸`,  `걹`,  `걺`,  `걻`,  `걼`,  `걽`,  `걾`,  `걿`,
  `！`,  `＂`,  `＃`,  `＄`,  `％`,  `＆`,  `＇`,  `（`,  `）`,  `＊`,  `＋`,  `，`,  `－`,  `．`,  `／`,  `０`,  `１`,  `２`,  `３`,  `４`,  `５`,  `６`,  `７`,  `８`,  `９`,  `：`,  `；`,  `＜`,  `＝`,  `＞`,  `？`,  `＠`,  `Ａ`,  `Ｂ`,  `Ｃ`,  `Ｄ`,  `Ｅ`,  `Ｆ`,  `Ｇ`,  `Ｈ`,  `Ｉ`,  `Ｊ`,  `Ｋ`,  `Ｌ`,  `Ｍ`,  `Ｎ`,  `Ｏ`,  `Ｐ`,  `Ｑ`,  `Ｒ`,  `Ｓ`,  `Ｔ`,  `Ｕ`,  `Ｖ`,  `Ｗ`,  `Ｘ`,  `Ｙ`,  `Ｚ`,  `［`,  `＼`,  `］`,  `＾`,  `＿`,  `｀`,  `ａ`,  `ｂ`,  `ｃ`,  `ｄ`,  `ｅ`,  `ｆ`,  `ｇ`,  `ｈ`,  `ｉ`,  `ｊ`,  `ｋ`,  `ｌ`,  `ｍ`,  `ｎ`,  `ｏ`,  `ｐ`,  `ｑ`,  `ｒ`,  `ｓ`,  `ｔ`,  `ｕ`,  `ｖ`,  `ｗ`,  `ｘ`,  `ｙ`,  `ｚ`,  `｛`,  `｜`,  `｝`,  `～`,  `｡`,  `｢`,  `｣`,  `､`,  `･`,  `ｦ`,  `ｧ`,  `ｨ`,  `ｩ`,  `ｪ`,  `ｫ`,  `ｬ`,  `ｭ`,  `ｮ`,  `ｯ`,  `ｰ`,  `ｱ`,  `ｲ`,  `ｳ`,  `ｴ`,  `ｵ`,  `ｶ`,  `ｷ`,  `ｸ`,  `ｹ`,  `ｺ`,  `ｻ`,  `ｼ`,  `ｽ`,  `ｾ`,  `ｿ`,  `ﾀ`,  `ﾁ`,  `ﾂ`,
  `Ο`, `ὐ`, `χ`, `ὶ`,  `τ`, `α`, `ὐ`, `τ`, `ὰ`,  `π`, `α`, `ρ`, `ί`, `σ`, `τ`, `α`, `τ`, `α`, `ί`,  `μ`, `ο`, `ι`,  `γ`, `ι`, `γ`, `ν`, `ώ`, `σ`, `κ`, `ε`, `ι`, `ν`, `,`,  `ὦ`,  `ἄ`, `ν`, `δ`, `ρ`, `ε`, `ς`,  `᾿`, `Α`, `θ`, `η`, `ν`, `α`, `ῖ`, `ο`, `ι`, `,`, 
  `ὅ`, `τ`, `α`, `ν`,  `τ`, `᾿`,  `ε`, `ἰ`, `ς`,  `τ`, `ὰ`,  `π`, `ρ`, `ά`, `γ`, `μ`, `α`, `τ`, `α`,  `ἀ`, `π`, `ο`, `β`, `λ`, `έ`, `ψ`, `ω`,  `κ`, `α`, `ὶ`,  `ὅ`, `τ`, `α`, `ν`,  `π`, `ρ`, `ὸ`, `ς`,  `τ`, `ο`, `ὺ`, `ς`, 
  `λ`, `ό`, `γ`, `ο`, `υ`, `ς`,  `ο`, `ὓ`, `ς`,  `ἀ`, `κ`, `ο`, `ύ`, `ω`, `·`,  `τ`, `ο`, `ὺ`, `ς`,  `μ`, `ὲ`, `ν`,  `γ`, `ὰ`, `ρ`,  `λ`, `ό`, `γ`, `ο`, `υ`, `ς`,  `π`, `ε`, `ρ`, `ὶ`,  `τ`, `ο`, `ῦ`, 
  `τ`, `ι`, `μ`, `ω`, `ρ`, `ή`, `σ`, `α`, `σ`, `θ`, `α`, `ι`,  `Φ`, `ί`, `λ`, `ι`, `π`, `π`, `ο`, `ν`,  `ὁ`, `ρ`, `ῶ`,  `γ`, `ι`, `γ`, `ν`, `ο`, `μ`, `έ`, `ν`, `ο`, `υ`, `ς`, `,`,  `τ`, `ὰ`,  `δ`, `ὲ`,  `π`, `ρ`, `ά`, `γ`, `μ`, `α`, `τ`, `᾿`,  
  `ε`, `ἰ`, `ς`,  `τ`, `ο`, `ῦ`, `τ`, `ο`,  `π`, `ρ`, `ο`, `ή`, `κ`, `ο`, `ν`, `τ`, `α`, `,`,   `ὥ`, `σ`, `θ`, `᾿`,  `ὅ`, `π`, `ω`, `ς`,  `μ`, `ὴ`,  `π`, `ε`, `ι`, `σ`, `ό`, `μ`, `ε`, `θ`, `᾿`,  `α`, `ὐ`, `τ`, `ο`, `ὶ`, 
  `π`, `ρ`, `ό`, `τ`, `ε`, `ρ`, `ο`, `ν`,  `κ`, `α`, `κ`, `ῶ`, `ς`,  `σ`, `κ`, `έ`, `ψ`, `α`, `σ`, `θ`, `α`, `ι`,  `δ`, `έ`, `ο`, `ν`, `.`,  `ο`, `ὐ`, `δ`, `έ`, `ν`,  `ο`, `ὖ`, `ν`,  `ἄ`, `λ`, `λ`, `ο`,  `μ`, `ο`, `ι`,  `δ`, `ο`, `κ`, `ο`, `ῦ`, `σ`, `ι`, `ν`, 
  `ο`, `ἱ`,  `τ`, `ὰ`,  `τ`, `ο`, `ι`, `α`, `ῦ`, `τ`, `α`,  `λ`, `έ`, `γ`, `ο`, `ν`, `τ`, `ε`, `ς`,  `ἢ`,  `τ`, `ὴ`, `ν`,  `ὑ`, `π`, `ό`, `θ`, `ε`, `σ`, `ι`, `ν`, `,`,  `π`, `ε`, `ρ`, `ὶ`,  `ἧ`, `ς`,  `β`, `ο`, `υ`, `λ`, `ε`, `ύ`, `ε`, `σ`, `θ`, `α`, `ι`, `,`, 
  `ο`, `ὐ`, `χ`, `ὶ`,  `τ`, `ὴ`, `ν`,  `ο`, `ὖ`, `σ`, `α`, `ν`,  `π`, `α`, `ρ`, `ι`, `σ`, `τ`, `ά`, `ν`, `τ`, `ε`, `ς`,  `ὑ`, `μ`, `ῖ`, `ν`,  `ἁ`, `μ`, `α`, `ρ`, `τ`, `ά`, `ν`, `ε`, `ι`, `ν`, `.`,  `ἐ`, `γ`, `ὼ`,  `δ`, `έ`, `,`,  `ὅ`, `τ`, `ι`,  `μ`, `έ`, `ν`, 
  `π`, `ο`, `τ`, `᾿`,  `ἐ`, `ξ`, `ῆ`, `ν`,  `τ`, `ῇ`,  `π`, `ό`, `λ`, `ε`, `ι`,  `κ`, `α`, `ὶ`,  `τ`, `ὰ`,  `α`, `ὑ`, `τ`, `ῆ`, `ς`,  `ἔ`, `χ`, `ε`, `ι`, `ν`,  `ἀ`, `σ`, `φ`, `α`, `λ`, `ῶ`, `ς`,  `κ`, `α`, `ὶ`,  `Φ`, `ί`, `λ`, `ι`, `π`, `π`, `ο`, `ν`, 
  `τ`, `ι`, `μ`, `ω`, `ρ`, `ή`, `σ`, `α`, `σ`, `θ`, `α`, `ι`, `,`,  `κ`, `α`, `ὶ`,  `μ`, `ά`, `λ`, `᾿`,  `ἀ`, `κ`, `ρ`, `ι`, `β`, `ῶ`, `ς`,  `ο`, `ἶ`, `δ`, `α`, `·`,  `ἐ`, `π`, `᾿`,  `ἐ`, `μ`, `ο`, `ῦ`,  `γ`, `ά`, `ρ`, `,`,  `ο`, `ὐ`,  `π`, `ά`, `λ`, `α`, `ι`, 
  `γ`, `έ`, `γ`, `ο`, `ν`, `ε`, `ν`,  `τ`, `α`, `ῦ`, `τ`, `᾿`,  `ἀ`, `μ`, `φ`, `ό`, `τ`, `ε`, `ρ`, `α`, `·`,  `ν`, `ῦ`, `ν`,  `μ`, `έ`, `ν`, `τ`, `ο`, `ι`,  `π`, `έ`, `π`, `ε`, `ι`, `σ`, `μ`, `α`, `ι`,  `τ`, `ο`, `ῦ`, `θ`, `᾿`,  `ἱ`, `κ`, `α`, `ν`, `ὸ`, `ν`, 
  `π`, `ρ`, `ο`, `λ`, `α`, `β`, `ε`, `ῖ`, `ν`,  `ἡ`, `μ`, `ῖ`, `ν`,  `ε`, `ἶ`, `ν`, `α`, `ι`,  `τ`, `ὴ`, `ν`,  `π`, `ρ`, `ώ`, `τ`, `η`, `ν`, `,`,  `ὅ`, `π`, `ω`, `ς`,  `τ`, `ο`, `ὺ`, `ς`,  `σ`, `υ`, `μ`, `μ`, `ά`, `χ`, `ο`, `υ`, `ς`, 
  `σ`, `ώ`, `σ`, `ο`, `μ`, `ε`, `ν`, `.`,  `ἐ`, `ὰ`, `ν`,  `γ`, `ὰ`, `ρ`,  `τ`, `ο`, `ῦ`, `τ`, `ο`,  `β`, `ε`, `β`, `α`, `ί`, `ω`, `ς`,  `ὑ`, `π`, `ά`, `ρ`, `ξ`, `ῃ`, `,`,  `τ`, `ό`, `τ`, `ε`,  `κ`, `α`, `ὶ`,  `π`, `ε`, `ρ`, `ὶ`,  `τ`, `ο`, `ῦ`, 
  `τ`, `ί`, `ν`, `α`,  `τ`, `ι`, `μ`, `ω`, `ρ`, `ή`, `σ`, `ε`, `τ`, `α`, `ί`,  `τ`, `ι`, `ς`,  `κ`, `α`, `ὶ`,  `ὃ`, `ν`,  `τ`, `ρ`, `ό`, `π`, `ο`, `ν`,  `ἐ`, `ξ`, `έ`, `σ`, `τ`, `α`, `ι`,  `σ`, `κ`, `ο`, `π`, `ε`, `ῖ`, `ν`, `·`,  `π`, `ρ`, `ὶ`, `ν`,  `δ`, `ὲ`, 
  `τ`, `ὴ`, `ν`,  `ἀ`, `ρ`, `χ`, `ὴ`, `ν`,  `ὀ`, `ρ`, `θ`, `ῶ`, `ς`,  `ὑ`, `π`, `ο`, `θ`, `έ`, `σ`, `θ`, `α`, `ι`, `,`,  `μ`, `ά`, `τ`, `α`, `ι`, `ο`, `ν`,  `ἡ`, `γ`, `ο`, `ῦ`, `μ`, `α`, `ι`,  `π`, `ε`, `ρ`, `ὶ`,  `τ`, `ῆ`, `ς`, 
  `τ`, `ε`, `λ`, `ε`, `υ`, `τ`, `ῆ`, `ς`,  `ὁ`, `ν`, `τ`, `ι`, `ν`, `ο`, `ῦ`, `ν`,  `π`, `ο`, `ι`, `ε`, `ῖ`, `σ`, `θ`, `α`, `ι`,  `λ`, `ό`, `γ`, `ο`, `ν`, `.`,
  `გ`, `თ`, `ხ`, `ო`, `ვ`, `თ`,  `ა`, `ხ`, `ლ`, `ა`, `ვ`, `ე`,  `გ`, `ა`, `ი`, `ა`, `რ`, `ო`, `თ`,  `რ`, `ე`, `გ`, `ი`, `ს`, `ტ`, `რ`, `ა`, `ც`, `ი`, `ა`,  `U`, `n`, `i`, `c`, `o`, `d`, `e`, `-`, `ი`, `ს`,  `მ`, `ე`, `ა`, `თ`, `ე`,  `ს`, `ა`, `ე`, `რ`, `თ`, `ა`, `შ`, `ო`, `რ`, `ი`, `ს`, `ო`, 
  `კ`, `ო`, `ნ`, `ფ`, `ე`, `რ`, `ე`, `ნ`, `ც`, `ი`, `ა`, `ზ`, `ე`,  `დ`, `ა`, `ს`, `ა`, `ს`, `წ`, `რ`, `ე`, `ბ`, `ა`, `დ`, `,`,  `რ`, `ო`, `მ`, `ე`, `ლ`, `ი`, `ც`,  `გ`, `ა`, `ი`, `მ`, `ა`, `რ`, `თ`, `ე`, `ბ`, `ა`,  `1`, `0`, `-`, `1`, `2`,  `მ`, `ა`, `რ`, `ტ`, `ს`, `,`, 
  `ქ`, `.`,  `მ`, `ა`, `ი`, `ნ`, `ც`, `შ`, `ი`, `,`,  `გ`, `ე`, `რ`, `მ`, `ა`, `ნ`, `ი`, `ა`, `შ`, `ი`, `.`,  `კ`, `ო`, `ნ`, `ფ`, `ე`, `რ`, `ე`, `ნ`, `ც`, `ი`, `ა`,  `შ`, `ე`, `ჰ`, `კ`, `რ`, `ე`, `ბ`, `ს`,  `ე`, `რ`, `თ`, `ა`, `დ`,  `მ`, `ს`, `ო`, `ფ`, `ლ`, `ი`, `ო`, `ს`, 
  `ე`, `ქ`, `ს`, `პ`, `ე`, `რ`, `ტ`, `ე`, `ბ`, `ს`,  `ი`, `ს`, `ე`, `თ`,  `დ`, `ა`, `რ`, `გ`, `ე`, `ბ`, `შ`, `ი`,  `რ`, `ო`, `გ`, `ო`, `რ`, `ი`, `ც`, `ა`, `ა`,  `ი`, `ნ`, `ტ`, `ე`, `რ`, `ნ`, `ე`, `ტ`, `ი`,  `დ`, `ა`,  `U`, `n`, `i`, `c`, `o`, `d`, `e`, `-`, `ი`, `,`, 
  `ი`, `ნ`, `ტ`, `ე`, `რ`, `ნ`, `ა`, `ც`, `ი`, `ო`, `ნ`, `ა`, `ლ`, `ი`, `ზ`, `ა`, `ც`, `ი`, `ა`,  `დ`, `ა`,  `ლ`, `ო`, `კ`, `ა`, `ლ`, `ი`, `ზ`, `ა`, `ც`, `ი`, `ა`, `,`,  `U`, `n`, `i`, `c`, `o`, `d`, `e`, `-`, `ი`, `ს`,  `გ`, `ა`, `მ`, `ო`, `ყ`, `ე`, `ნ`, `ე`, `ბ`, `ა`, 
  `ო`, `პ`, `ე`, `რ`, `ა`, `ც`, `ი`, `უ`, `ლ`,  `ს`, `ი`, `ს`, `ტ`, `ე`, `მ`, `ე`, `ბ`, `ს`, `ა`, `,`,  `დ`, `ა`,  `გ`, `ა`, `მ`, `ო`, `ყ`, `ე`, `ნ`, `ე`, `ბ`, `ი`, `თ`,  `პ`, `რ`, `ო`, `გ`, `რ`, `ა`, `მ`, `ე`, `ბ`, `შ`, `ი`, `,`,  `შ`, `რ`, `ი`, `ფ`, `ტ`, `ე`, `ბ`, `შ`, `ი`, `,`, 
  `ტ`, `ე`, `ქ`, `ს`, `ტ`, `ე`, `ბ`, `ი`, `ს`,  `დ`, `ა`, `მ`, `უ`, `შ`, `ა`, `ვ`, `ე`, `ბ`, `ა`, `ს`, `ა`,  `დ`, `ა`,  `მ`, `რ`, `ა`, `ვ`, `ა`, `ლ`, `ე`, `ნ`, `ო`, `ვ`, `ა`, `ნ`,  `კ`, `ო`, `მ`, `პ`, `ი`, `უ`, `ტ`, `ე`, `რ`, `უ`, `ლ`,  `ს`, `ი`, `ს`, `ტ`, `ე`, `მ`, `ე`, `ბ`, `შ`, `ი`, `.`,
	]
)
